library verilog;
use verilog.vl_types.all;
entity Packet_sv_unit is
end Packet_sv_unit;

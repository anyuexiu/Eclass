library verilog;
use verilog.vl_types.all;
entity data_defs_v_unit is
end data_defs_v_unit;

interface TA_Probe_io(
	//Fetch In
	input logic enable_updatePC_in,
	input logic enable_fetch_in,
	input logic [15:0] taddr_in,
	input logic br_taken_in,
	//Fetch Out
	input logic [15:0] pc2cmp,
	input logic [15:0] npc2cmp,
	input logic IMem_rd2cmp,
	//Decode In
	input logic [15:0] IMem_dout_in,
	input logic [15:0] npc_in_in,
//	input logic [2:0] psr_in,
	input logic enable_decode_in,
	//Decode Out
	input logic [15:0] IR2cmp,
	input logic [15:0] npc_out2cmp,
	input logic [5:0] E_control2cmp,
	input logic [1:0] W_control2cmp,
	input logic Mem_control2cmp,
	//Execute in
	input logic enable_execute_in,
	input logic [5:0] E_control_in,
	input logic bypass_alu_1_in,
	input logic bypass_alu_2_in,
	input logic bypass_mem_1_in,
	input logic bypass_mem_2_in,
	input logic [15:0] IR_in,
	input logic [15:0] ex_npc_in,
	input logic  Mem_control_in,
	//input logic [1:0] W_control_in,
	input logic [15:0] VSR1_in,
	input logic [15:0] VSR2_in,
	input logic [15:0] mem_bypass_in,
	input logic [15:0] aluout_prev_in,
	//Execute Out
	input logic [1:0] W_Control_out2cmp,
	input logic  Mem_Control_out2cmp,
	input logic [15:0] aluout2cmp,
	input logic [2:0] dr2cmp,
	input logic [2:0] sr12cmp,
	input logic [2:0] sr22cmp,
	//input logic alucarry2cmp,
	input logic [2:0] NZP2cmp,
	input logic [15:0] IR_Exec2cmp,
	input logic [15:0] M_Data2cmp,
	input logic [15:0] imm52cmp,
	input logic [15:0] offset62cmp, 
	input logic [15:0] offset92cmp, 
	input logic [15:0] offset112cmp,
	
	//Writeback inputs
	input logic enable_wb_in,
	input logic [1:0] W_Control_wb_in,
	input logic [15:0] pcout_wb_in,
	input logic [15:0] memout_wb_in,
	input logic [2:0] dr_wb_in,
	input logic [2:0] sr1_wb_in,
	input logic [2:0] sr2_wb_in,
	input logic [15:0] npc_wb_in,
	input logic [15:0] aluout_wb_in,
	input logic [15:0] ram_wb_in[0:7],
	//Writeback outputs
	input logic [15:0] VSR12cmp,
	input logic [15:0] VSR22cmp,
	input logic [2:0] psr2cmp,
	//Controller inputs
	input logic complete_data_in,
	input logic complete_instr_in,
	input logic [15:0] IR_ctrl_in,
	input logic [15:0] IR_Exec_in,
	input logic [2:0] NZP_in,
	input logic [2:0] psr_in,
	//Controller outputs
	input logic enable_updatePC2cmp,
	input logic enable_fetch2cmp,
	input logic enable_decode2cmp,
	input logic enable_execute2cmp,
	input logic enable_writeback2cmp,
	input logic bypass_alu_12cmp,
	input logic bypass_alu_22cmp,
	input logic bypass_mem_12cmp,
	input logic bypass_mem_22cmp,
	input logic [1:0] mem_state2cmp,
	input logic br_taken2cmp,
	//Memaccess Inputs
	input logic [1:0] mem_state_in,
	input logic  M_control_in,
	input logic [15:0] M_Data_in,	
	input logic [15:0] M_Addr_in,
	input logic [15:0] Data_dout_in,
	//Memaccess Outputs
	input logic [15:0] Data_addr2cmp,
  	input logic [15:0] Data_din2cmp,
  	input logic Data_rd2cmp,
  	input logic [15:0] memout2cmp
	//Cache Inputs
	//input logic dmac,
	//input logic rd,
	//input logic [15:0] addr,
	//input logic [15:0] din,
	//input logic rrdy,
	//input logic rdrdy,
	//input logic wacpt,
	//input logic miss_in,
	//input logic [3:0] state_in,
	//input logic [1:0] count_in,
	//input logic [63:0] blockdata_in,
	//input logic valid_in,
	//input logic [15:0] offdata_in,
	//input logic [15:0] validarr_in,
	//input logic [73:0] memdata_in,
	//Cache Outpus
	//input logic [15:0] dout,
	//input logic complete,
	//input logic rrqst,
	//input logic rdacpt,
	//input logic wrqst,
	//input logic [15:0] offdata_out,
	//input logic miss_out,
	//input logic [3:0] state_out,
	//input logic [1:0] count_out,
	//input logic [63:0] blockdata_out,
	//input logic valid_out,
	//input logic [15:0] validarr_out,
	//input logic ramrd_out,
	//input logic [63:0] blkreg_out
);
endinterface


library verilog;
use verilog.vl_types.all;
entity Execute_test_top is
    generic(
        simulation_cycle: integer := 10
    );
end Execute_test_top;

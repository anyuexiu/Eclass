library verilog;
use verilog.vl_types.all;
entity Execute_test is
    generic(
        reg_wd          : integer := 32
    );
end Execute_test;

library verilog;
use verilog.vl_types.all;
entity LC3_io is
    port(
        clock           : in     vl_logic
    );
end LC3_io;

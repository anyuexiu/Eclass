library verilog;
use verilog.vl_types.all;
entity Execute_if_sv_unit is
end Execute_if_sv_unit;

library verilog;
use verilog.vl_types.all;
entity LC3_test is
    generic(
        reg_wd          : integer := 16
    );
end LC3_test;
